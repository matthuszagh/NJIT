PACKAGE n_bit_int IS
    SUBTYPE S9  IS INTEGER RANGE -2**8  TO 2**8-1;
    SUBTYPE S11 IS INTEGER RANGE -2**10 TO 2**10-1;
    SUBTYPE S15 IS INTEGER RANGE -2**14 TO 2**14-1;
    SUBTYPE S16 IS INTEGER RANGE -2**15 TO 2**15-1;
    SUBTYPE S22 IS INTEGER RANGE -2**21 TO 2**21-1;
    SUBTYPE S30 IS INTEGER RANGE -2**29 TO 2**29-1;
    SUBTYPE S32 IS INTEGER RANGE -2**31 TO 2**31-1;
END PACKAGE;
