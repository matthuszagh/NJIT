-- fft8.vhd
--
-- A 8-length FFT using the Cooley-Tukey algorithm.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

USE work.n_bit_int.ALL;
--------------------------------------------------------------------------------
ENTITY fft8 IS
    GENERIC (LENGTH : INTEGER := 8;    -- Filter length.
             STAGES : INTEGER := 3     -- M=lg(LENGTH)
    );
    PORT (clk     : IN  STD_LOGIC;
          reset   : IN  STD_LOGIC;
          x_in    : IN  S10;
          X_r_out : OUT A0_7S10;
          X_i_out : OUT A0_7S10
    );
END ENTITY fft8;
--------------------------------------------------------------------------------
ARCHITECTURE fpga OF fft8 IS

    TYPE CONST_ARR IS ARRAY (0 TO STAGES) OF A0_2S17;
    TYPE A0_M_A0_7S10 IS ARRAY (0 TO STAGES) OF A0_7S10;

    CONSTANT W : CONST_ARR := 
            (( 32768,  32768,  32768),  -- 1
             ( 23170,      0,  46340),  -- cos( pi/4) - isin( pi/4)
             (     0, -32768,  32768),  -- -i
             (-23170,      0, -46340)); -- cos(3pi/4) - isin(3pi/4)

    SIGNAL count : INTEGER RANGE -1 TO LENGTH-1 := LENGTH-1;
    SIGNAL xmr   : A0_M_A0_7S10 := (OTHERS => (OTHERS => 0)); -- Array at stage M - reals
    SIGNAL xmi   : A0_M_A0_7S10 := (OTHERS => (OTHERS => 0)); -- Array at stage M - imaginaries

    COMPONENT butterfly IS
        PORT (clk    : IN  STD_LOGIC;
              reset  : IN  STD_LOGIC;
              in1_r  : IN  S10;
              in1_i  : IN  S10;
              in2_r  : IN  S10;
              in2_i  : IN  S10;
              tw_r   : IN  S17;
              tw_rpi : IN  S17;
              tw_rmi : IN  S17;
              out1_r : OUT S10;
              out1_i : OUT S10;
              out2_r : OUT S10;
              out2_i : OUT S10
        );
    END COMPONENT butterfly;

BEGIN

    load_x: PROCESS (clk, reset) IS
    BEGIN
        IF reset='1' THEN
            --xmr <= (OTHERS => (OTHERS => 0));
            --xmi <= (OTHERS => (OTHERS => 0));
            count  <= LENGTH-1;
        ELSIF rising_edge(clk) THEN
            IF count >= 0 THEN
                xmr(0)(LENGTH-1) <= x_in;
                FOR i IN LENGTH-1 DOWNTO 1 LOOP
                    xmr(0)(i-1) <= xmr(0)(i);
                END LOOP;
                count <= count-1;
            END IF;
        END IF;
    END PROCESS load_x;

    -- Perform butterfly computations in every stage.
    stage: FOR i IN 0 TO STAGES-1 GENERATE
        substage: FOR j IN 0 TO LENGTH/2-1 GENERATE
            SIGNAL vec_index : UNSIGNED(STAGES-1 DOWNTO 0) := (OTHERS => '0');
            CONSTANT index : INTEGER RANGE 0 TO LENGTH-1
                    := TO_INTEGER(insert_pad_bit(reverse_vector(delete_bit(vec_index, STAGES-1-i)+j), STAGES-1-i));
            CONSTANT inc : INTEGER RANGE 1 TO LENGTH/2 := LENGTH/(2**(i+1));
            CONSTANT w_inc : UNSIGNED(1 DOWNTO 0) := TO_UNSIGNED(inc*j, 2);
        BEGIN
            butterfly_comp: butterfly
                PORT MAP (clk    => clk,
                          reset  => reset,
                          in1_r  => xmr(i)(index),
                          in1_i  => xmi(i)(index),
                          in2_r  => xmr(i)(index+inc),
                          in2_i  => xmi(i)(index+inc),
                          tw_r   => W(TO_INTEGER(w_inc))(0),
                          tw_rpi => W(TO_INTEGER(w_inc))(1),
                          tw_rmi => W(TO_INTEGER(w_inc))(2),
                          out1_r => xmr(i+1)(index),
                          out1_i => xmi(i+1)(index),
                          out2_r => xmr(i+1)(index+inc),
                          out2_i => xmi(i+1)(index+inc));
        END GENERATE substage;
    END GENERATE stage;

    -- Map internal data to output.
    output: FOR i IN 0 TO LENGTH-1 GENERATE
        SIGNAL vec_index : UNSIGNED(STAGES-1 DOWNTO 0) := (OTHERS => '0');
        CONSTANT index : INTEGER RANGE 0 TO LENGTH-1
                := TO_INTEGER(reverse_vector(vec_index+i));
    BEGIN
        X_r_out(i)            <= xmr(STAGES)(index);
        X_i_out(i)            <= xmi(STAGES)(index);
    END GENERATE output;

END ARCHITECTURE fpga;
